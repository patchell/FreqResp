N 7
R 1 6 3000.0
R 2 6 4700.0
A 6 1 6 2 0.15
R 0 1 250000.0
R 1 3 68000.0
R 3 5 68000.0
C 5 2 0.00001
C 3 6 0.0000001
C 1 4 0.000000001
C 4 5 0.000000001
R 4 6 400000.0
I 0
O 2
G 6
S 1.0 7 20

