N 3
R 0 1 1.0
C 1 2 1.0
I 0
O 1
G 2
S 0.1 2 10

