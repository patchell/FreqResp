N 8
R 0 1 10000.0
R 1 2 10000.0
A 3 1 7 2 100.0
R 2 7 100.0
R 0 3 10000.0
C 3 7 0.0000001

R 2 4 10000.0
R 4 5 10000.0
A 6 4 7 5 100.0
R 5 7 100.0
R 2 6 10000.0
C 6 7 0.00004

I 0
O 5
G 7
S 0.1 5 20

