N 5
R 0 1 10000.0
R 1 2 10000.0
A 3 1 4 2 100.0
R 2 4 100.0
R 0 3 10000.0
C 3 4 0.0000001
I 0
O 2
G 4
S 1.0 4 20

