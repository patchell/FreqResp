N 3
R 0 2 1.0
R 1 2 2.0
A 2 0 2 1 1.0
I 0
O 1
G 2
S 1.0 2 5

