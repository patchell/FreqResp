N 4
R 0 1 1.0
L 1 2 1.0
C 2 3 1.0
I 0
O 2
G 3
S 0.1 2 30
