R 0 1 20000.0
R 1 2 20000.0
C 1 4 0.0000001
C 0 3 0.000000001
C 3 2 0.000000001
R 3 4 400.0
N 5
I 0
O 2
S 100.0 4 10
G 4

